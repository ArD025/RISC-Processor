module processor(clk1, clk2);  // only the inputs are clk1 and clk2
input clk1, clk2;  // two phase clocks
reg [31:0] PC, IF_ID_IR, IF_ID_NPC;  // registers of stage 1
reg [31:0] ID_EX_NPC, ID_EX_IR, ID_EX_A, ID_EX_B, ID_EX_Imm;  // registers of stage 2
reg [2:0] ID_EX_type, EX_MEM_type, MEM_WB_type;  // type of instructions like R-R R-Imm
reg [31:0] EX_MEM_ALUOUT, EX_MEM_IR, EX_MEM_B;  // register of stage 3
reg EX_MEM_cond;  // condition for branch
reg [31:0] MEM_WB_IR, MEM_WB_ALUOUT, MEM_WB_LMD;
reg [31:0] regfile[31:0];  // register bank of 32 register with each register having data of 32 bits
reg [31:0] mem[1023:0];  // memory file of 1204 words with each word of 32 bits
reg HALTED;  // when halt is executed then HALTED is set to 1 when it reaches the stage WB 
reg TAKEN_BRANCH; // when TAKEN_BRANCH is set to 1 then all the instructions entered the pipeline are disabled or they write nothing on registers and memory

// Below are the operations(func) specifies by 6 bit opcode in IR
parameter ADD=6'b000000, SUB=6'b000001, AND=6'b000010, OR=6'b000011, SLT=6'b000100, MUL=6'b000101, HLT=6'b111111, LW=6'b001000, SW=6'b001001;
parameter ADDI=6'b001010, SUBI=6'b001011, SLTI=6'b001100, BNEQZ=6'b001101, BEQZ=6'b001110; 

// Below are the types of instructions given by the opcode
parameter RR_ALU=3'b000, RM_ALU=3'b001, LOAD=3'b010, STORE=3'b011, BRANCH=3'b100, HALT=3'b101;

// lets write the code of IF stage which works on posedge of clk1
always@ (posedge clk1)
begin
if(HALTED==0)  // if HALTED==1 then the whole program is skipped out
begin
if(((EX_MEM_IR[31:26]==BEQZ) && EX_MEM_cond==1)|| ((EX_MEM_IR[31:26]==BNEQZ) && EX_MEM_cond==))
begin
IF_ID_IR <= #2 mem[EX_MEM_ALUOUT];
TAKEN_BRANCH <= #2 1'b1;
IF_ID_NPC <= #2 EX_MEM_ALUOUT+1;
PC <= #2 EX_MEM_ALUOUT;
end
else
begin
IF_ID_IR <= #2 mem[PC];
IF_ID_NPC <= #2 PC+1;
PC <= #2 PC+1;
end
end
end

// lets write the code of ID stage which works on posedge of clk2
always@ (posedge clk2)
begin
if(HALTED==0)
begin
if(IF_ID_IR[25:21]==5'b00000)
begin
ID_EX_A <= 0;
end
else
begin
ID_EX_A <= #2 regfile[IF_ID_IR[25:21]];  // rs
end
if(IF_ID_IR[20:16]==5'b00000)
begin
ID_EX_B <= 0;
end
else
begin
ID_EX_B <= #2 regfile[IF_ID_IR[20:16]];  // rt
end
ID_EX_IR <= #2 IF_ID_IR;
ID_EX_NPC <= #2 IF_ID_NPC;
ID_EX_Imm <= #2 {{16{IF_ID_IR[15]}},IF_ID_IR[15:0]};  // sign extend Imm
end

// Now lets see what type of instruction is given to us
case(IF_ID_IR[31:26])
ADD, SUB, AND, OR, MUL, SLT: ID_EX_type <= #2 RR_ALU;
ADDI, SUBI, SLTI :           ID_EX_type <= #2 RM_ALU;
LW:                          ID_EX_type <= #2 LOAD;
SW:                          ID_EX_type <= #2 STORE;
BNEQZ, BEQZ:                 ID_EX_type <= #2 BRANCH;
HLT:                         ID_EX_type <= #2 HALT;
default:                     ID_EX_type <= #2 HALT;  // invalid opcode
endcase
end

// Lets write the code of EX stage which works on posedge clk2
always@ (posedge clk1)
begin
if(HALTED==0)
begin
EX_MEM_IR <= #2 ID_EX_IR;
EX_MEM_type <= #2 ID_EX_type;
TAKEN_BRANCH <= #2 1'b0;  // TAKEN_BRANCH is initialized to 0
case(ID_EX_type)
RR_ALU: begin
case(ID_EX_IR[31:26])
ADD: 	 EX_MEM_ALUOUT <= #2 ID_EX_A + ID_EX_B;
SUB: 	 EX_MEM_ALUOUT <= #2 ID_EX_A - ID_EX_B;
AND: 	 EX_MEM_ALUOUT <= #2 ID_EX_A & ID_EX_B;
OR:  	 EX_MEM_ALUOUT <= #2 ID_EX_A | ID_EX_B;
MUL: 	 EX_MEM_ALUOUT <= #2 ID_EX_A * ID_EX_B;
SLT: 	 EX_MEM_ALUOUT <= #2 ID_EX_A < ID_EX_B;
default: EX_MEM_ALUOUT <= #2 32'bxxxxxxxx;
endcase
end
RM_ALU: begin
case(ID_EX_IR[31:26])
ADDI:  	 EX_MEM_ALUOUT <= #2 ID_EX_A + ID_EX_Imm;
SUBI: 	 EX_MEM_ALUOUT <= #2 ID_EX_A - ID_EX_Imm;
SLTI: 	 EX_MEM_ALUOUT <= #2 ID_EX_A < ID_EX_Imm;
default: EX_MEM_ALUOUT <= #2 32'bxxxxxxxx;
endcase
end
LOAD, STORE: begin
EX_MEM_ALUOUT <= #2 ID_EX_A + ID_EX_Imm;
EX_MEM_B <= #2 ID_EX_B;
end
BRANCH: begin
EX_MEM_ALUOUT <= #2 ID_EX_NPC + ID_EX_Imm;
EX_MEM_cond <= #2 (ID_EX_A==0);
BEQZ: EX_MEM_cond <= #2 (ID_EX_A == 0);
BNEQZ: EX_MEM_cond <= #2 (ID_EX_A != 0);
end
endcase
end
end

// Lets write a code of MEM stage which works on posedge of clk2
always@ (posedge clk2)
begin
if(HALTED==0)
begin
MEM_WB_type <= #2 EX_MEM_type;
MEM_WB_IR <= #2 EX_MEM_IR;
case(EX_MEM_type)
RR_ALU, RM_ALU: MEM_WB_ALUOUT <= #2 EX_MEM_ALUOUT;
LOAD: MEM_WB_LMD <= #2 mem[EX_MEM_ALUOUT];
STORE: begin
if(TAKEN_BRANCH==0)  // Disable writing on register and memory
mem[EX_MEM_ALUOUT] <= #2 EX_MEM_B;
end
endcase
end
end

// Lets write code of WB stage which works on posedge clk1
always@ (posedge clk1)
begin
if(TAKEN_BRANCH==0)
begin
case(MEM_WB_type)
RR_ALU: regfile[MEM_WB_IR[15:11]] <= #2 MEM_WB_ALUOUT;
RM_ALU: regfile[MEM_WB_IR[20:16]] <= #2 MEM_WB_ALUOUT;
LOAD: regfile[MEM_WB_IR[20:16]] <= #2 MEM_WB_LMD;
HALT: HALTED <= #2 1'b1;
endcase
end
end
endmodule
