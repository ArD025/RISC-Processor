
module testbench;
reg clk1, clk2;
integer k;
processor DUT(clk1, clk2);
initial
begin
clk1=0;
forever       // generating of two phase clock pulses
begin
#5 clk1=1;
#5 clk1=0;
#10 clk1=0;
end
end
initial
begin
clk2=0;
forever
begin
#15 clk2=1;
#5 clk2=0;
end
end
initial
begin
for(k=0; k<32; k=k+1)
DUT.regfile[k]=k;
end
initial
begin
DUT.mem[0]=32'h28010078;
DUT.mem[1]=32'h0c631800;
DUT.mem[2]=32'h20220000;
DUT.mem[3]=32'h0c631800;
DUT.mem[4]=32'h2842002d;
DUT.mem[5]=32'h0c631800;
DUT.mem[6]=32'h24220001;
DUT.mem[7]=32'hfc000000;
DUT.mem[120]=85;
end
initial
begin
DUT.PC=0;
DUT.HALTED=0;
DUT.TAKEN_BRANCH=0;
$dumpfile("processor.vcd");
$dumpvars(0, testbench);
#500 $monitor("mem[120] = %1d \nmem[121] = %1d", DUT.mem[120], DUT.mem[121]);
#10 $finish;
end
endmodule
